/**
*******************************************************************************
* @file    mod_main.sv
* @author  Victor Hugo Becerril Bueno
* @email   vhugobeb@gmail.com
* @brief   This is a simple example of a D type flip flop as the
*          main module of the project.
*******************************************************************************
* @Description
* This is a simple example of a D-type flip flop as the main module of the
* project. Where the data type that goes through the circuit is composed of a
* tag and a data, this data type is declared in the definitions.svh file.
*
*******************************************************************************
*/

/*****************************************************************************/
/*          START OF INCLUDES                                                */
/*****************************************************************************/
`include "definitions.svh"
/*****************************************************************************/
/*          END OF INCLUDES                                                  */
/*****************************************************************************/

/*****************************************************************************/
/*          START OF MAIN MODULE                                             */
/*****************************************************************************/
module mod_main(
    // Inputs
    input          i_clk,             // Enable Signal
    input            i_E,             // Enable Signal
    input  Bus_t     i_D,             // Data Input
    // Outputs
    output Bus_t     o_Q,             // Data Output
    output Bus_t    o_nQ              // Output data denied
);

    /*************************************************************************/
    /*          START OF REGISTERS                                           */
    /*************************************************************************/
    /*************************************************************************/
    /*          END OF REGISTERS                                             */
    /*************************************************************************/

    /*************************************************************************/
    /*          START OF WIRES                                               */
    /*************************************************************************/
    /*************************************************************************/
    /*          END OF WIRES                                                 */
    /*************************************************************************/

    /*************************************************************************/
    /*          START OF BITS                                                */
    /*************************************************************************/
    /*************************************************************************/
    /*          END OF BITS                                                  */
    /*************************************************************************/

    /*************************************************************************/
    /*          START OF SEQUENTIAL PROCESS                                  */
    /*************************************************************************/
    always_ff @( posedge i_clk ) begin : D_Type_Flip_Flop
        if ( i_E ) begin
            o_Q  <= i_D;
        end
        else begin
            o_Q  <= 12'b0;
        end
    end : D_Type_Flip_Flop
    /*************************************************************************/
    /*          END OF SEQUENTIAL PROCESS                                    */
    /*************************************************************************/

    /*************************************************************************/
    /*          START OF COMBINATORIAL PROCESS                               */
    /*************************************************************************/
    assign o_nQ = ~o_Q;
    /*************************************************************************/
    /*          END OF COMBINATORIAL PROCESS                                 */
    /*************************************************************************/

endmodule
/*****************************************************************************/
/*          END OF MAIN MODULE                                               */
/*****************************************************************************/
