/**
******************************************************************************
* @file    definitions.svh
* @author  Victor Hugo Becerril Bueno
* @email   vhugobeb@gmail.com
* @brief   Definition of the project
******************************************************************************
* @Description
* This is an example of header file for declareate datatypes and macros
*
******************************************************************************
*/

`ifndef DEFINITIONS_SVH_
`define DEFINITIONS_SVH_

/*****************************************************************************/
/*          START OF DEFINES                                                 */
/*****************************************************************************/
/*****************************************************************************/
/*          END OF DEFINES                                                   */
/*****************************************************************************/

/*****************************************************************************/
/*           START OF MACROS                                                 */
/*****************************************************************************/
/*****************************************************************************/
/*           END OF MACROS                                                   */
/*****************************************************************************/

/*****************************************************************************/
/*          START OF DATATYPES                                               */
/*****************************************************************************/
/*
* @brief:        Bus_t structure definition
* @description:  This contains a Tag and Data value
*/
typedef struct packed {
    logic [ 3 : 0 ] Tag;
    logic [ 7 : 0 ] Data;
} Bus_t;
/*****************************************************************************/
/*          END OF DATATYPES                                                 */
/*****************************************************************************/
`endif  /* DEFINITIONS_SVH_ */
